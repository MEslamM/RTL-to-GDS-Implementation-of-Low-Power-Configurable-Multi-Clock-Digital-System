`timescale 1ns/1ns  
module Full_System_TB ();

/////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////declare testbench signals////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////

reg              i_clk_ref = 1 ;  
reg              i_clk_UART = 1 ;  
reg				 i_rx_in ;
reg              i_rst ; 
wire        	 o_tx_out ;
wire        	 o_parr_err ;
wire        	 o_fram_err ;

integer 		 i ;
/////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////clocks///////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////

parameter ref_clk_period = 20 ; //50Mhz
parameter UART_clk_period = 200 ; //5Mhz

/////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////test cases//////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////

//Writing In Reg commands (1st TEST CASE)
reg [0:10] Writing_Reg_command = 11'b0_01010101_0_1 ; //'haa+even_parity (mirror)
reg [0:10] address_Reg_command = 11'b0_00000101_0_1 ; //Address = 5
reg [0:10] data_Reg_command = 11'b0_00000101_0_1 ; //data = 5

//Reading From Reg Commands (2nd TEST CASE)
reg [0:10] Reading_Reg_command = 11'b0_11011101_0_1 ; //'hbb+even_parity (read address 5) (mirror)

//Testing ALU with operands (3rd TEST CASE)
reg [0:10] ALU_OPERANDS_command = 11'b0_00110011_0_1 ; //'hcc+even_parity (mirror)
reg [0:10] OP_A_Value_command = 11'b0_11000000_0_1 ; //Value =3 (mirror)
reg [0:10] OP_B_Value_command = 11'b0_11000000_0_1 ; //Value =3 (mirror)
reg [0:10] Function_Value_command = 11'b0_0000000_0_1 ; //Adder (mirror)

/////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////// Clock Generator////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////

always #(ref_clk_period/2) i_clk_ref = ~i_clk_ref  ;  
always #(UART_clk_period/2) i_clk_UART = ~i_clk_UART  ; 

/////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////Module declaration //////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////

Final_system DUT0(
 .RST_N(i_rst),
 .UART_CLK(i_clk_UART),
 .REF_CLK(i_clk_ref),
 .UART_RX_IN(i_rx_in),
 .UART_TX_O(o_tx_out),
 .parity_error(o_parr_err),
 .framing_error(o_fram_err)
);

/////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////initial block////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////

initial begin 
i_rst=0;
i_rx_in=1;
#900
i_rst=1;
#300
/////////////////////////////////////////////////////////////////////////////////////////

//Testing Writing in Reg case 
for ( i = 0; i < 11; i=i+1) begin
i_rx_in=Writing_Reg_command[i];
#1600;
end

#800
for ( i = 0; i < 11; i=i+1) begin
i_rx_in=address_Reg_command[i];
#1600;
end

#800
for ( i = 0; i < 11; i=i+1) begin
i_rx_in=data_Reg_command[i];
#1600;
end

#1000
/////////////////////////////////////////////////////////////////////////////////////////

//Testing Reading from Reg case 
for ( i = 0; i < 11; i=i+1) begin
i_rx_in=Reading_Reg_command[i];
#1600;
end

#800
for ( i = 0; i < 11; i=i+1) begin
i_rx_in=address_Reg_command[i];
#1600;
end

#62000
/////////////////////////////////////////////////////////////////////////////////////////

//Tetsing ALU With operands
for ( i = 0; i < 11; i=i+1) begin
i_rx_in=ALU_OPERANDS_command[i];
#1600;
end

#800
for ( i = 0; i < 11; i=i+1) begin
i_rx_in=OP_A_Value_command[i];
#1600;
end

#800
for ( i = 0; i < 11; i=i+1) begin
i_rx_in=OP_B_Value_command[i];
#1600;
end

#800
for ( i = 0; i < 11; i=i+1) begin
i_rx_in=Function_Value_command[i];
#1600;
end
/////////////////////////////////////////////////////////////////////////////////////////

#62000


$stop;
end


endmodule